`include "types/decoupled.sv"
