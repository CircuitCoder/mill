`include "utils/mem_arbiter.sv"

module instr_fetch;
endmodule
