`ifndef __EXECUTE_SV__
`define __EXECUTE_SV__

`include "types.sv"

`endif // __EXECUTE_SV__
